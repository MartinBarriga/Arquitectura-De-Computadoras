library ieee;
use ieee.std_logic_1164.all;
library lattice;
use lattice.component.all;

entity adder